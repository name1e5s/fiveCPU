`timescale 1ns / 1ps
module alu_alpha(
        input   clk,
        input   rst,
        
        input   [31:0] a,
        input   [31:0] b,
        output   [63:0] c
    );
    
    
endmodule
